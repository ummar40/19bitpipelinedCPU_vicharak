//Also we've a parameter.v module which defines many parametes as:
`define ART 5'd0
`define LOG 5'd1
`define JMP 5'd2
`define BQE 5'd3
`define BNE 5'd4
`define CALL 5'd5
`define RET 5'd6
`define LD 5'd7
`define ST 5'd8
`define CRY 5'd9
`define IMM 5'd10

`define ADD 5'd0
`define SUB 5'd1
`define MUL 5'd2
`define DIV 5'd3
`define INC 5'd4
`define DEC 5'd5
`define AND 5'd6
`define OR 5'd7
`define XOR 5'd8
`define NOT 5'd9
`define ENCRY 5'd10
`define DECRY 5'd11
`define IMMED 5'd12